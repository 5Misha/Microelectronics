
`timescale 1ns / 1ps

module tb_counter_2bit;

logic clk_t, _rst_t;
logic [7:0] Q_t;

top DUT ( .clk(clk_t), ._rst(_rst_t), .Q(Q_t) );

// Генератор тактового сигнала
initial begin
    clk_t = 0;
    for (int i = 0; i < 50; i++) begin
        #5 clk_t = ~clk_t;
    end
end

// Тестовые воздействия
initial begin
    // Инициализация
    _rst_t = 0;
    #20 _rst_t = 1;
    $display("Time\tTens\tUnits");
    $monitor("%0d\t%0d\t%0d", $time, Q_t[7:4], Q_t[3:0]);

    // Сброс
    #120 _rst_t = 0;
    #10 _rst_t = 1;
    #40;

end

endmodule